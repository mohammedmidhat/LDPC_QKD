//////////////////////////////////////////////////////////////////////////////////
// Company:         MIT Quantum Photonics Group
// Author:        	Mohammed Al Ai Baky
// 
// Create Date:     6/6/2018 
// Design Name:     LDPC_decoder_Frolov_1024_0.5
// Module Name:     top 
// Project Name:    LDPC_decoder_Frolov_1024_0.5
// Target Devices:  VC707 Virtex-7 FPGA
// Tool versions:   Vivado 2017.4
// Description:     top module for the LDPC decoder
//
// Dependencies: 	decoder_2048_1024.v
//					clock_divider.v
//
// Revision: 
// Revision 0.0
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module top#(parameter max_iter = 30, parameter log2max_iter = 5, parameter INT = 8, parameter FRAC = 8, parameter deg_v = 7, parameter deg_c = 10,
				parameter circ = 128, parameter log2circ = 8, parameter n = 2048)(
	input clk_p,
	input clk_n,
	input rst,
	output success,
	output [log2max_iter-1:0] iterations
	);

IBUFDS #(
    .DIFF_TERM("FALSE"), // Differential Termination
    .IBUF_LOW_PWR("TRUE"), // Low power="TRUE", Highest perforrmance="FALSE"
    .IOSTANDARD("DEFAULT") // Specify the input I/O standard
    ) IBUFDS_inst (
    .O(clk_in), // Buffer output
    .I(clk_p), // Diff_p buffer input (connect directly to top-level port)
    .IB(clk_n) // Diff_n buffer input (connect directly to top-level port)
    );

clock_divider clock_divider_inst(
	.clk_in(clk_in),
	.clk_out(clk_out)
	);

decoder decoder_inst(
	.clk(clk_out),
	.rst(rst),
	.data(2048'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000100000000000000000000010000000000100000000000000000001000000000000000000001000000000000000000000000000000100000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000010000010000000000000000000000000000000000000000000000001000001000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000001000001000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000001000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000100000000000000000100000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000010000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000001000000000100000001000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000010000000000000000000000010000000000010000000000000001000000000000000000000000),
	.success(success),
	.iterations(iterationso)
	);

endmodule
