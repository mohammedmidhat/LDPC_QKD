module decoder#(parameter n = 204, parameter m = 102, parameter log2n = 8, parameter log2m = 7, parameter max_iter = 30, parameter log2max_iter = 5,
				parameter INT = 8, parameter FRAC = 8, parameter deg_v = 3, parameter deg_c = 6, parameter log2deg_v = 2, parameter log2deg_c = 3)(
	input clk,
	input rst,
	output success,
	output [log2max_iter-1:0] iterations
	);

wire [n*deg_v*log2m-1:0] v_neighbor;
wire [m*deg_c*log2n-1:0] c_neighbor;
wire [m*deg_c*log2deg_v-1:0] neighbor_index_to_var;	// specifies the neighboring index of a check to a var
													// e.g. ch2 is the 1st neighbor check in its 3rd var neighbor
wire [n*deg_v*log2deg_c-1:0] neighbor_index_to_ch;	// specifies the neighboring index of a var to a check
													// e.g. var2 is the 1st neighbor check in its 3rd check neighbor
assign v_neighbor = 4284'b110010010100000000111001000101001100000011010010010011111001011011010101010111010001110000010111010001011010100111000101011011011111001110100000110011101100100001010110001101101011100011110100111001111111001001010101100011000001001001110110001101010000101001110101101001100000001101001000010100000100110100100001110101010101000100100111001110010100111000111010110101010011010111000101110000011011100101000000110101010010100100111001100101001101110101011001011001010001000010101001111101101010111100010111011100101100100000100011011011001000011101001010110100010001101001001001110110011000000111101011110110111101001010110010100000000110000111101001000000010000000011000110011101000100100111001110001101011011000010101010000110011100110100011010110111000001100000000111011011000000000100101100001010101011100000101000101001001110000110110001100110110101110011001110001001001011011111100111100001000010001010000100010001011101001111110001111000000011000001001110101011100010110111000111101011100000001110011111000011110001000100100000011001100110100010101011010101010101111010011001100000101110011001000110001011010010111101000000101000000110110000001100101101101100001101001010001000001101101001101010111010001011100100000101010110001011110001101010010000111011100101001000110000101010110000101000100011101100100011111100010110000100010111000100110011010110100111010001111000100110110011000100000011010010011100101101110001010011100001000101011100000101000101111100000001011001110011010010101001100110000100110101100001110010010110100011110000101111010100001010001010100001111100000101101000100110100010001111010011011000010101000010100101101100010111110100001100110011001010010000011110100111001100001010100000010011000011011011110010111100011110010100110111010101010101011000001001110011111101100010011100001011010010100111111101111001010000101100000111011000010111000001100010101000001100010010100111110010010010001111000110110010001011100001010111110100011101101110101010101110000000110110110000001010011100001000010000001111000110000010011101110010011010101111110011000111100011000101101010000010011010000011100010110100100000100010101101010000001010100001101010001001000001000110001000000011101010000011001101111001010110101000111001010011101011110110110111000010100000100011000000011000011001110011000011001101000110010111010101011110110011000000100001001100000101010110000101101011011101010001101011100001010010111000010000001001110011000011011011100001010010101011011010000010010000010011011100001110010100001100010011110010001010010000101001010000011001101101010111011000101100011010111000010001110001101100011001000001001100100000000110110010001110101011011101000011000001010101110010101111100010100010101011001001001001001111011000111100001000110010110100011100011010011000011001111011011010101110000111011101010010010101111011101110111110111101101110100001100011111101111001101101100101101010101110111010100101111100111110000001010111101010110101101100000000101110101110000001100101010111011100111010101100001110010100110001100111110100110001101110000010000111010100111100010000101101100100010011001100010111100110101101100101001100001000100010000101001010111001101101101001011110110001000110111000111011100111001101001110101100001000110001111010110100011110111001011001001001001011001010010110000100110110011000110000000010000011011101000010110011000110100000101100000100011110011100100111000011100111010101000001011100111100010101001100101001011001100100100001000100100101001001010001000110010011100010001010001011101110000110101001010010110000100010110000110000000111001100110011010110011000100100000100001110000000100001110000001011001101100010100000110011110010000101111011010011000001000000010010111010101110100101001011000000110011110100110101010010010110100000010010010000110000101100111100001111011000101001101100110110001001010100100100111000001111100101100101011000010100100110101001001011001011000111100011000000110001011111100101100010110010110000111101010010100010001110100010010100001100110110001111000001101011010110001100011101101110100010010010010100010100001000100101001011000100111111011110000001001100100010011001001110100011011111001111110101100000100100010100110100100101001011110011000001000110011010110111011111101011010011010100100110101001010001;
assign c_neighbor = 4896'b010110001000110000110011101110000010001010101010010011000111100101100010011111010100001110010110010011101100110001001011101100110000100010010011010100001010101101001010011100010000110001111010001101001010001100001001110001110011101010001110010110111000110101001000011101000100101001111100001000101100100001001101011110000010110010001000010000010110101001000101011111100001000110100011010000110111010100111000101101010011010110010010010001001011011101010010110010000101101110100001001001000110111001010001100111100101100010111010000010111001010101100001101010010100111011000111010100101011010101001001100011000101011110011000001101111000111001011101101011110011000010110111001100100111111000001100100100100001011110101000010111011010011001000111101001000011011010111011000011001001101000111101110000000110001111000101010000101011110101010111100110100100110101111001000110011010101000000001011100110100001010000011000101101100000000111010101111000001110110001001000010011010111100011011101111100101010010111001011000101000011100001011101100100000000111001001010011011011100100001010110011000110010011000001000101111010001000011010110010100100100010110110001111011100001100101011011011010011001101111000000011011010010000000011100001100001111110010100001110110111110100100001011010100010100011000000000100001000100100011001011110100001101111001010000001001001000001010101011101100010010010010101000000011011100001000110100001000100101111000011001001110110011101010100100100010101000010101110001010110110111100001101101000000011010010111100010100011010100100111100110000010110010110101101000111101001111000100101100100110101001010100110001101101000000000100110100111000000101010001101010101011000010000011000101001010101111101111011010111001000100000101111100001010110000110101011011000001000000101010110101110100000110110101001001111111010100000101110100101100101110110100000000000100111011100000110110000110000100101110110000001101100011001001100100001110011110001110000011000010111110000011101100000000100010110011110000010001000001101100011011011000001001001101010010001011100010101000010101100010011111010010001010001101010110001001110110001100101111010001100001100111011010001011111011010110011000110101100001001011001110100100000100010010001010101110100001011010111101000111011011011110000001110110000010001111011001101000011100101000010111101101110001000011100100101011011011010010011100010000101010010000110100000110101100000010000010110000100011000111000011000010110100110110010110110001011001100001001100000111001101101000010011001110001001011100110100101010000011101110001011010100101000100011001111101011100100110010010001101101100010000001001011100000100101100000100011010011010010110011001001101011010110001000011111110011001001100011011101100000010101010110100000001100111001000111000111100010010101101110000011001110101000110111100001001000000110010010001010010011111010010110111100001100110100000100101110001101111001111001100011100001111101110110001001110111000000010100111101101010011011101010010101010010111010101000110101100000111100111110010101110111101000001111001100100110111110010110001101010000001001011110111001000101000101000110010011101111111000110001100101000110000101111110010000110011100010110100111000100110010100100000000011110001111011001011011011000100111101111010000111110011011000111011010000100101101011111110000111001111110011001100110110001100101100101110001100110101111000101001010000001000001011100100100010010011101010010101000101100101001101011100001111011000100000011101100000100101010101010000110001010110011000111111011110000100010011111000100100101110111001101011100010000110100011110010101011010000000010111101001000100100100101110010000001001101011001010001000010101011110101010100101001110100100001110000111001100010001100110000000010010110001001010010111000000111111100000110001110010110101000100100111011000010100101001110001000001101000000101011011001000111110100010000010100110000110010101111000001000110110100011110100110010111111010011111010010100010011100010110011100110001010001001101011000100010101101011000000101101110010000000111100101100100011011001110101000110100010011001001001010001001111110001010010111001111101000011111011000000110001100011100011001010000010001110100111010001100100011010000011110110111110001011001001011001011000100010100110011010110010010010011010111001100000110000100101010101110011001110011011101000010000100011010010010111001000010100111001001000000101101101100101101010100111000001011011111000001110011110110101100111000010001000001000101001011001101000010011011101101101001010101001110000010111100111010100011111001100010111111001101101000100100101010100111111000110000100110111111100011111011100000001100010010000010101101010110100001000101000100010000010110100001111101011111100011110011011100110000011001011000111000110110100101100101001100011101101101001000110101010011100011100101011010100000110000111;
assign neighbor_index_to_var = 1224'b000001011010000001011010000001011010000001011010000001011010000001011010000001011010000001011010000001011010000001011010000001011010000001011010000001011010000001011010000001011010000001011010000001011010000001011010000001011010000001011010000001011010000001011010000001011010000001011010000001011010000001011010000001011010000001011010000001011010000001011010000001011010000001011010000001011010000001011010000001011010000001011010000001011010000001011010000001011010000001011010000001011010000001011010000001011010000001011010000001011010000001011010000001011010000001011010000001011010000001011010000001011010000001011010000001011010000001011010000001011010000001011010000001011010000001011010000001011010000001011010000001011010000001011010000001011010000001011010000001011010000001011010000001011010000001011010000001011010000001011010000001011010000001011010000001011010000001011010000001011010000001011010000001011010000001011010000001011010000001011010000001011010000001011010000001011010000001011010000001011010000001011010000001011010000001011010000001011010000001011010000001011010000001011010000001011010000001011010000001011010000001011010000001011010000001011010000001011010000001011010000001011010000001011010;
assign neighbor_index_to_ch = 1836'b001011101001011101001011101001011101001011101001011101001011101001011101001011101001011101001011101001011101001011101001011101001011101001011101001011101001011101001011101001011101001011101001011101001011101001011101001011101001011101001011101001011101001011101001011101001011101001011101001011101001011101001011101001011101001011101001011101001011101001011101001011101001011101001011101001011101001011101001011101001011101001011101001011101001011101001011101001011101001011101001011101001011101001011101001011101001011101001011101001011101001011101001011101001011101001011101001011101001011101001011101001011101001011101001011101001011101001011101001011101001011101001011101001011101001011101001011101001011101001011101001011101001011101001011101001011101001011101001011101001011101001011101001011101001011101001011101001011101001011101001011101001011101001011101001011101001011101001011101001011101001011101001011101000010100000010100000010100000010100000010100000010100000010100000010100000010100000010100000010100000010100000010100000010100000010100000010100000010100000010100000010100000010100000010100000010100000010100000010100000010100000010100000010100000010100000010100000010100000010100000010100000010100000010100000010100000010100000010100000010100000010100000010100000010100000010100000010100000010100000010100000010100000010100000010100000010100000010100000010100000010100000010100000010100000010100000010100000010100000010100000010100000010100000010100000010100000010100000010100000010100000010100000010100000010100000010100000010100000010100000010100000010100000010100000010100000010100000010100000010100000010100000010100000010100000010100000010100000010100000010100000010100000010100000010100000010100000010100000010100000010100000010100000010100000010100000010100000010100000010100000010100000010100000010100000010100;

reg [n*deg_v*(INT+FRAC)-1:0] v_msg;
reg [m*deg_c*(INT+FRAC)-1:0] c_msg;
wire [INT+FRAC-1:0] LLR = 16'b1010101011001011;
reg [n*(INT+FRAC)-1:0] LLRs;

wire [n-1:0] data = 12'b100101010101;
reg [n-1:0] dec_cw;
reg [2:0] FSM;
reg non_zero_syn;

reg success_dec;
assign success = success_dec;

reg [log2max_iter-1:0] iter_num;
assign iterations = iter_num;
reg [log2n-1:0] data_iter;
reg [log2m-1:0] check_iter;


wire [log2deg_v-1:0] neighbor_index_to_var_5;
wire [log2deg_v-1:0] neighbor_index_to_var_4;
wire [log2deg_v-1:0] neighbor_index_to_var_3;
wire [log2deg_v-1:0] neighbor_index_to_var_2;
wire [log2deg_v-1:0] neighbor_index_to_var_1;
wire [log2deg_v-1:0] neighbor_index_to_var_0;

wire [log2n-1:0] vn_5_ind;
wire [log2n-1:0] vn_4_ind;
wire [log2n-1:0] vn_3_ind;
wire [log2n-1:0] vn_2_ind;
wire [log2n-1:0] vn_1_ind;
wire [log2n-1:0] vn_0_ind;

assign neighbor_index_to_var_5 = neighbor_index_to_var[((check_iter+1)*deg_c)*log2deg_v-1 -: log2deg_v];
assign neighbor_index_to_var_4 = neighbor_index_to_var[((check_iter+1)*deg_c-1)*log2deg_v-1 -: log2deg_v];
assign neighbor_index_to_var_3 = neighbor_index_to_var[((check_iter+1)*deg_c-2)*log2deg_v-1 -: log2deg_v];
assign neighbor_index_to_var_2 = neighbor_index_to_var[((check_iter+1)*deg_c-3)*log2deg_v-1 -: log2deg_v];
assign neighbor_index_to_var_1 = neighbor_index_to_var[((check_iter+1)*deg_c-4)*log2deg_v-1 -: log2deg_v];
assign neighbor_index_to_var_0 = neighbor_index_to_var[((check_iter+1)*deg_c-5)*log2deg_v-1 -: log2deg_v];

assign vn_5_ind = c_neighbor[((check_iter+1)*deg_c)*log2n-1 -: log2n];
assign vn_4_ind = c_neighbor[((check_iter+1)*deg_c-1)*log2n-1 -: log2n];
assign vn_3_ind = c_neighbor[((check_iter+1)*deg_c-2)*log2n-1 -: log2n];
assign vn_2_ind = c_neighbor[((check_iter+1)*deg_c-3)*log2n-1 -: log2n];
assign vn_1_ind = c_neighbor[((check_iter+1)*deg_c-4)*log2n-1 -: log2n];
assign vn_0_ind = c_neighbor[((check_iter+1)*deg_c-5)*log2n-1 -: log2n];

reg [INT+FRAC-1:0] vn_cn_msgs_0_5;
reg [INT+FRAC-1:0] vn_cn_msgs_0_4;
reg [INT+FRAC-1:0] vn_cn_msgs_0_3;
reg [INT+FRAC-1:0] vn_cn_msgs_0_2;
reg [INT+FRAC-1:0] vn_cn_msgs_0_1;
reg [INT+FRAC-1:0] vn_cn_msgs_0_0;

reg [INT+FRAC-1:0] cn_vn_msgs_2;
reg [INT+FRAC-1:0] cn_vn_msgs_1;
reg [INT+FRAC-1:0] cn_vn_msgs_0;

wire [INT+FRAC-1:0] cn_vn_msgs_0_0;
wire [INT+FRAC-1:0] cn_vn_msgs_0_1;
wire [INT+FRAC-1:0] cn_vn_msgs_0_2;
wire [INT+FRAC-1:0] cn_vn_msgs_0_3;
wire [INT+FRAC-1:0] cn_vn_msgs_0_4;
wire [INT+FRAC-1:0] cn_vn_msgs_0_5;

wire [INT+FRAC-1:0] vn_out_1;
wire [INT+FRAC-1:0] vn_out_2;
wire [INT+FRAC-1:0] vn_out_3;
wire [INT+FRAC-1:0] belief_out;

reg bit_0_in;
reg bit_1_in;
reg bit_2_in;
reg bit_3_in;
reg bit_4_in;
reg bit_5_in;
wire syn_res;


cn cn_0_inst (
	.msg_in_1(vn_cn_msgs_0_0),
	.msg_in_2(vn_cn_msgs_0_1),
	.msg_in_3(vn_cn_msgs_0_2),
	.msg_in_4(vn_cn_msgs_0_3),
	.msg_in_5(vn_cn_msgs_0_4),
	.msg_in_6(vn_cn_msgs_0_5),
	.msg_out_1(cn_vn_msgs_0_0),
	.msg_out_2(cn_vn_msgs_0_1),
	.msg_out_3(cn_vn_msgs_0_2),
	.msg_out_4(cn_vn_msgs_0_3),
	.msg_out_5(cn_vn_msgs_0_4),
	.msg_out_6(cn_vn_msgs_0_5)
	);

vr vn_0_inst (
	.ch_msg_0(cn_vn_msgs_0),
	.ch_msg_1(cn_vn_msgs_1),
	.ch_msg_2(cn_vn_msgs_2),
	.vr_msg_0(vn_out_1),
	.vr_msg_1(vn_out_2),
	.vr_msg_2(vn_out_3),
	.belief(belief_out)
	);

syn	syn_0_inst (
	.bit_0(bit_0_in),
	.bit_1(bit_1_in),
	.bit_2(bit_2_in),
	.bit_3(bit_3_in),
	.bit_4(bit_4_in),
	.bit_5(bit_5_in),
	.result(syn_res)
	);


always @(posedge clk or posedge rst) begin
	if (rst) begin
		FSM <= 0;
		success_dec <= 0;
		data_iter <= 1;
		check_iter <= 1;
		iter_num <= 0;
		dec_cw <= data;
		non_zero_syn <= 0;
	end

	else if (FSM == 0) begin
		if (data_iter < n+1) begin
			LLRs[data_iter*(INT+FRAC)-1 -: INT+FRAC] <= data[data_iter-1]*LLR;
		
			v_msg[data_iter*deg_v*(INT+FRAC)-1 -: INT+FRAC] <= data[data_iter-1]*LLR;
			v_msg[(data_iter*deg_v-1)*(INT+FRAC)-1 -: INT+FRAC] <= data[data_iter-1]*LLR;
			v_msg[(data_iter*deg_v-2)*(INT+FRAC)-1 -: INT+FRAC] <= data[data_iter-1]*LLR;

			data_iter <= data_iter + 1;
		end
		
		if(data_iter == n+1)begin
			data_iter <= 1;
			FSM <= 1;

			vn_cn_msgs_0_5 <= v_msg[((c_neighbor[(deg_c)*log2n-1 -: log2n])*deg_v-neighbor_index_to_var[(deg_c)*log2deg_v-1 -: log2deg_v])*(INT+FRAC)-1 -: INT+FRAC];
			vn_cn_msgs_0_4 <= v_msg[((c_neighbor[(deg_c-1)*log2n-1 -: log2n])*deg_v-neighbor_index_to_var[(deg_c-1)*log2deg_v-1 -: log2deg_v])*(INT+FRAC)-1 -: INT+FRAC];
			vn_cn_msgs_0_3 <= v_msg[((c_neighbor[(deg_c-2)*log2n-1 -: log2n])*deg_v-neighbor_index_to_var[(deg_c-2)*log2deg_v-1 -: log2deg_v])*(INT+FRAC)-1 -: INT+FRAC];
			vn_cn_msgs_0_2 <= v_msg[((c_neighbor[(deg_c-3)*log2n-1 -: log2n])*deg_v-neighbor_index_to_var[(deg_c-3)*log2deg_v-1 -: log2deg_v])*(INT+FRAC)-1 -: INT+FRAC];
			vn_cn_msgs_0_1 <= v_msg[((c_neighbor[(deg_c-4)*log2n-1 -: log2n])*deg_v-neighbor_index_to_var[(deg_c-4)*log2deg_v-1 -: log2deg_v])*(INT+FRAC)-1 -: INT+FRAC];
			vn_cn_msgs_0_0 <= v_msg[((c_neighbor[(deg_c-5)*log2n-1 -: log2n])*deg_v-neighbor_index_to_var[(deg_c-5)*log2deg_v-1 -: log2deg_v])*(INT+FRAC)-1 -: INT+FRAC];

			bit_5_in <= dec_cw[c_neighbor[(deg_c)*log2n-1 -: log2n]];
			bit_4_in <= dec_cw[c_neighbor[(deg_c-1)*log2n-1 -: log2n]];
			bit_3_in <= dec_cw[c_neighbor[(deg_c-2)*log2n-1 -: log2n]];
			bit_2_in <= dec_cw[c_neighbor[(deg_c-3)*log2n-1 -: log2n]];
			bit_1_in <= dec_cw[c_neighbor[(deg_c-4)*log2n-1 -: log2n]];
			bit_0_in <= dec_cw[c_neighbor[(deg_c-5)*log2n-1 -: log2n]];
		end
	end

	else if (FSM == 1) begin
		if (check_iter < m+1) begin
			check_iter <= check_iter + 1;

			c_msg[check_iter*deg_c*(INT+FRAC)-1 -: INT+FRAC] <= cn_vn_msgs_0_5;
			c_msg[(check_iter*deg_c-1)*(INT+FRAC)-1 -: INT+FRAC] <= cn_vn_msgs_0_4;
			c_msg[(check_iter*deg_c-2)*(INT+FRAC)-1 -: INT+FRAC] <= cn_vn_msgs_0_3;
			c_msg[(check_iter*deg_c-3)*(INT+FRAC)-1 -: INT+FRAC] <= cn_vn_msgs_0_2;
			c_msg[(check_iter*deg_c-4)*(INT+FRAC)-1 -: INT+FRAC] <= cn_vn_msgs_0_1;
			c_msg[(check_iter*deg_c-5)*(INT+FRAC)-1 -: INT+FRAC] <= cn_vn_msgs_0_0;

			if(syn_res) begin
				non_zero_syn <= 1;
			end
		end

		if (check_iter < m) begin
			vn_cn_msgs_0_5 <= v_msg[(vn_5_ind*deg_v-neighbor_index_to_var_5)*(INT+FRAC)-1 -: INT+FRAC];
			vn_cn_msgs_0_4 <= v_msg[(vn_4_ind*deg_v-neighbor_index_to_var_4)*(INT+FRAC)-1 -: INT+FRAC];
			vn_cn_msgs_0_3 <= v_msg[(vn_3_ind*deg_v-neighbor_index_to_var_3)*(INT+FRAC)-1 -: INT+FRAC];
			vn_cn_msgs_0_2 <= v_msg[(vn_2_ind*deg_v-neighbor_index_to_var_2)*(INT+FRAC)-1 -: INT+FRAC];
			vn_cn_msgs_0_1 <= v_msg[(vn_1_ind*deg_v-neighbor_index_to_var_1)*(INT+FRAC)-1 -: INT+FRAC];
			vn_cn_msgs_0_0 <= v_msg[(vn_0_ind*deg_v-neighbor_index_to_var_0)*(INT+FRAC)-1 -: INT+FRAC];

			bit_5_in <= dec_cw[vn_5_ind];
			bit_4_in <= dec_cw[vn_4_ind];
			bit_3_in <= dec_cw[vn_3_ind];
			bit_2_in <= dec_cw[vn_2_ind];
			bit_1_in <= dec_cw[vn_1_ind];
			bit_0_in <= dec_cw[vn_0_ind];
		end

		if(check_iter == m+1)begin
			check_iter <= 1;
			FSM <= 2;

			cn_vn_msgs_2 <= c_msg[((v_neighbor[(deg_v)*log2m-1 -: log2m])*deg_c-neighbor_index_to_ch[(deg_v)*log2deg_c-1 -: log2deg_c])*(INT+FRAC)-1 -: INT+FRAC];
			cn_vn_msgs_1 <= c_msg[((v_neighbor[(deg_v-1)*log2m-1 -: log2m])*deg_c-neighbor_index_to_ch[(deg_v-1)*log2deg_c-1 -: log2deg_c])*(INT+FRAC)-1 -: INT+FRAC];
			cn_vn_msgs_0 <= c_msg[((v_neighbor[(deg_v-2)*log2m-1 -: log2m])*deg_c-neighbor_index_to_ch[(deg_v-2)*log2deg_c-1 -: log2deg_c])*(INT+FRAC)-1 -: INT+FRAC];
		end
	end

	else if(FSM == 2) begin
		if(non_zero_syn) begin
			FSM <= 3;
			iter_num <= iter_num + 1;
		end else begin
			FSM <= 4;
		end
	end

	else if(FSM == 3) begin
		if(iter_num < max_iter) begin
			if (data_iter < n+1) begin
				data_iter <= data_iter + 1;

				v_msg[data_iter*deg_v*(INT+FRAC)-1 -: INT+FRAC] <= vn_out_3;
				v_msg[(data_iter*deg_v-1)*(INT+FRAC)-1 -: INT+FRAC] <= vn_out_2;
				v_msg[(data_iter*deg_v-2)*(INT+FRAC)-1 -: INT+FRAC] <= vn_out_1;

				dec_cw[data_iter] <= ~belief_out[INT+FRAC-1];
			end

			if (data_iter < n) begin
				cn_vn_msgs_2 <= c_msg[((v_neighbor[((data_iter+1)*deg_v)*log2m-1 -: log2m])*deg_c-neighbor_index_to_ch[((data_iter+1)*deg_v)*log2deg_c-1 -: log2deg_c])*(INT+FRAC)-1 -: INT+FRAC];
				cn_vn_msgs_1 <= c_msg[((v_neighbor[((data_iter+1)*deg_v-1)*log2m-1 -: log2m])*deg_c-neighbor_index_to_ch[((data_iter+1)*deg_v-1)*log2deg_c-1 -: log2deg_c])*(INT+FRAC)-1 -: INT+FRAC];
				cn_vn_msgs_0 <= c_msg[((v_neighbor[((data_iter+1)*deg_v-2)*log2m-1 -: log2m])*deg_c-neighbor_index_to_ch[((data_iter+1)*deg_v-2)*log2deg_c-1 -: log2deg_c])*(INT+FRAC)-1 -: INT+FRAC];
			end

			if (data_iter == n+1) begin
				data_iter <= 1;
				FSM <= 1;

				vn_cn_msgs_0_5 <= v_msg[((c_neighbor[(deg_c)*log2n-1 -: log2n])*deg_v-neighbor_index_to_var[(deg_c)*log2deg_v-1 -: log2deg_v])*(INT+FRAC)-1 -: INT+FRAC];
				vn_cn_msgs_0_4 <= v_msg[((c_neighbor[(deg_c-1)*log2n-1 -: log2n])*deg_v-neighbor_index_to_var[(deg_c-1)*log2deg_v-1 -: log2deg_v])*(INT+FRAC)-1 -: INT+FRAC];
				vn_cn_msgs_0_3 <= v_msg[((c_neighbor[(deg_c-2)*log2n-1 -: log2n])*deg_v-neighbor_index_to_var[(deg_c-2)*log2deg_v-1 -: log2deg_v])*(INT+FRAC)-1 -: INT+FRAC];
				vn_cn_msgs_0_2 <= v_msg[((c_neighbor[(deg_c-3)*log2n-1 -: log2n])*deg_v-neighbor_index_to_var[(deg_c-3)*log2deg_v-1 -: log2deg_v])*(INT+FRAC)-1 -: INT+FRAC];
				vn_cn_msgs_0_1 <= v_msg[((c_neighbor[(deg_c-4)*log2n-1 -: log2n])*deg_v-neighbor_index_to_var[(deg_c-4)*log2deg_v-1 -: log2deg_v])*(INT+FRAC)-1 -: INT+FRAC];
				vn_cn_msgs_0_0 <= v_msg[((c_neighbor[(deg_c-5)*log2n-1 -: log2n])*deg_v-neighbor_index_to_var[(deg_c-5)*log2deg_v-1 -: log2deg_v])*(INT+FRAC)-1 -: INT+FRAC];

				bit_5_in <= dec_cw[c_neighbor[(deg_c)*log2n-1 -: log2n]];
				bit_4_in <= dec_cw[c_neighbor[(deg_c-1)*log2n-1 -: log2n]];
				bit_3_in <= dec_cw[c_neighbor[(deg_c-2)*log2n-1 -: log2n]];
				bit_2_in <= dec_cw[c_neighbor[(deg_c-3)*log2n-1 -: log2n]];
				bit_1_in <= dec_cw[c_neighbor[(deg_c-4)*log2n-1 -: log2n]];
				bit_0_in <= dec_cw[c_neighbor[(deg_c-5)*log2n-1 -: log2n]];
			end
		end
	end

	else if(FSM == 4) begin
		success_dec <= 1;
	end
end

endmodule
